`include"gray_counter.v"
module tb_gray_counter(clk,rst,count);
reg clk,rst;
wire [2:0]
